--Michael Lange, 301580599; Trevor Ruttan, 301580889; Rohin Gill, 301582525;

library IEEE;
use ieee.std_logic_1164.all;

entity Part3 is 
	port (

			SW : in std_logic_vector(9 downto 0);
			HEX0, HEX1 : out std_logic_vector(6 downto 0)
			);
	end Part3;
	
architecture behavorial of Part3 is 
	begin
	end behavorial;