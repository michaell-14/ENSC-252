--------------------------------------
--Testbench tutorial
--Course: ENSC 252
--Original Creator: Anita Tino
--Edited: Sahaj Singh
---------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;

--declare a testbench. Testbench Entity is always empty
ENTITY oddCounter_tb IS
END oddCounter_tb;

ARCHITECTURE Behaviour of oddCounter_tb IS
	COMPONENT oddCounter IS --the component or DEVICE UNDER TEST (DUT) we would like to verify
	PORT(x1, x2, x3, x4 : IN STD_LOGIC;
			f : OUT STD_LOGIC);
	END COMPONENT;
	
	--signals used to connect above component to testbench
	--apply stimulus to input signals (seen below in stimulus process)
	--we view the output signals on the waveform, and verify that the DUT behaves as expected
	SIGNAL in1, in2, in3, in4, out_f : STD_LOGIC; 
	
	BEGIN
	
	DUT : oddCounter --declare the device under test (DUT) to be OddThing
	PORT MAP(x1 => in1, x2 => in2, x3 =>in3, x4 => in4, f => out_f); --map test signals to DUT
	
	stimulus : process
	BEGIN
		in1 <= '0'; --assign test stimulus "0000"
		in2 <= '0';
		in3 <= '0';
		in4 <= '0';
		--notice the space between "20 ns" 
		wait for 20 ns; --wait for data to propagate. See if expected output is generated by f in waveform
		
		in4 <= '1'; --assign test stimulus "0001"
		wait for 20 ns;

		in4 <= '0'; --assign test stimulus "0010"
		in3 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '0';
		in2 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '0';
		in2 <= '0';
		in1 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '0';
		in2 <= '1';	
		wait for 20 ns;

		in4 <= '1';
		wait for 20 ns;

		in4 <= '0';
		in3 <= '1';
		wait for 20 ns;

		in4 <= '1';
		wait for 100 ns;
		
		assert false;
		report "simulation ended" severity failure; --brute force quit so simulation does not run forever
		
		--Note: we can also use "assert" statements to create intelligent testbenches. EX:
		--wait for 20 ns;
		--assert f = '1';  
		--report "f is incorrect. Expected 1 when in1 = 0, in2 = ..." severity failure; 

		--report statements will be output to the Modelsim terminal window during simulation, which can help you 
		--pinpoint the issue in your waveform and design

		
	END process;
END Behaviour;
